module REG_FILE(
    input [4:0] read_reg_num1,
    input [4:0] read_reg_num2,
    input [4:0] write_reg,
    input [31:0] write_data,
    output reg [31:0] read_data1,
    output reg [31:0] read_data2,
    input regwrite,
    input clock,
    input reset
);

    reg [31:0] reg_memory [31:0];
    integer i;


    always @(posedge clock or posedge reset)
    begin
        if (reset) begin
            for (i = 0; i < 32; i = i + 1) begin
                reg_memory[i] <= 0;
            end
            read_data1 <= 0;
            read_data2 <= 0;
        end
        else begin
            if (regwrite && (write_reg != 5'b0)) begin
                reg_memory[write_reg] <= write_data;
            end

            read_data1 <= (read_reg_num1 == 5'b0) ? 32'h0 : reg_memory[read_reg_num1];
            read_data2 <= (read_reg_num2 == 5'b0) ? 32'h0 : reg_memory[read_reg_num2];
        end
    end


endmodule